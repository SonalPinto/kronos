// Copyright (c) 2020 Sonal Pinto
// SPDX-License-Identifier: Apache-2.0

/*
Kronos Hazard Control Unit

The HCU monitors for Register Read hazards at the Decode Stage
These hazards occur when a register is being read before it's
latest value is written back from the Write Back stage,
either as a result of a Direct Write or a Load

*/


module kronos_hcu 
    import kronos_types::*;
(
    input  logic        clk,
    input  logic        rstz,
    input  logic        flush,
    // Decoder inputs
    input  logic [4:0]  rs1,
    input  logic [4:0]  rs2,
    input  logic [4:0]  rd,
    input  logic        regrd_rs1_en,
    input  logic        regrd_rs2_en,
    input  logic        upgrade,
    // Write Back inputs
    input  logic [4:0]  regwr_sel,
    input  logic        downgrade,
    // Decoder Stall & forward status
    output logic        rs1_forward,
    output logic        rs2_forward,
    output logic        stall
);

/*
Register Pending Tracker
------------------------
In the Kronos pipeline, there are 2 stages ahead of the Decoder.

Hence, there can be a maximum of two pending writes to any register.

This is tracked as 2b shift register which shifts in a '1' to track
that a write is pending, and shifts out when it is written back.

This is representative of upgrading or downgrading the hazard level
on that register.

The LSB of this 2b hazard vector indicates the hazard status.

Controls,
Upgrade     : decode is ready to register for the next stage, and regwr_rd_en is valid
Downgrade   : write back is valid, i.e. regwr_en

Note,
1. This HCU design scales really well. For deeper levels of 
pending write-backs (downgrades), the hazard vector needs to be widened.
However, the stall condition only checks the LSB.

2. Register forwarding is possible when the hazard level is 1

This architecture can pretty much be used anywhere and at any stage if the IO is generalized

*/

logic [31:0][1:0] rpend;
logic rs1_stall, rs2_stall;

always_ff @(posedge clk or negedge rstz) begin
    if (~rstz) begin
        rpend <= '0;
    end
    else begin
        if (flush) begin
            rpend <= '0;
        end
        else if (upgrade && ~downgrade) begin
            // Decode ready. Upgrade register's hazard level
            rpend[rd] <= {rpend[rd][0], 1'b1};
        end
        else if (~upgrade && downgrade) begin
            // Register written back. Downgrade register's hazard level
            rpend[regwr_sel] <= {1'b0, rpend[regwr_sel][1]};
        end
        else if (upgrade && downgrade) begin
            // Hazard level remains the same if both decoder and write
            // back collide on the same register
            // Else, upgrade and downgrade specified registers
            if (rd != regwr_sel) begin
                rpend[rd] <= {rpend[rd][0], 1'b1};
                rpend[regwr_sel] <= {1'b0, rpend[regwr_sel][1]};
            end
        end
    end
end

// Detect register forwarding
assign rs1_forward = downgrade && rs1 == regwr_sel && rpend[rs1] == 2'b01;
assign rs2_forward = downgrade && rs2 == regwr_sel && rpend[rs2] == 2'b01;

// Stall conditions
assign rs1_stall = regrd_rs1_en && rpend[rs1][0] && ~rs1_forward;
assign rs2_stall = regrd_rs2_en && rpend[rs2][0] && ~rs2_forward;

// Stall if rs1 or rs2 is pending, and the register operands aren't being forwarded
assign stall = rs1_stall || rs2_stall;

endmodule